--------------------------------------------------------------------------------
--! @file top.vhd
--! @brief Toplevel module for TE0741-2C1.
--! @author Yuan Mei
--!
--! Target Devices: Kintex-7 XC7K160T-FFG676-2
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
LIBRARY UNISIM;
USE UNISIM.VComponents.ALL;

LIBRARY work;
USE work.utility.ALL;

ENTITY top IS
  GENERIC (
    ENABLE_DEBUG       : boolean := false;
    ENABLE_TEN_GIG_ETH : boolean := false
  );
  PORT (
    SYS_RST          : IN    std_logic;
    SYS_CLK_P        : IN    std_logic;
    SYS_CLK_N        : IN    std_logic;
    SGMIICLK_Q0_P    : IN    std_logic;  --! 125 MHz, for GTP/GTH/GTX
    SGMIICLK_Q0_N    : IN    std_logic;
    --
    LED8Bit          : OUT   std_logic_vector(7 DOWNTO 0);
    -- SFP
    SFP_TX_P         : OUT   std_logic;
    SFP_TX_N         : OUT   std_logic;
    SFP_RX_P         : IN    std_logic;
    SFP_RX_N         : IN    std_logic;
    SFP_LOS_LS       : IN    std_logic;
    SFP_TX_DISABLE_N : OUT   std_logic;
    -- MGT
    MGT_CLK3_P       : IN    std_logic;  --! 156.25 MHz, for GTX/10GbE
    MGT_CLK3_N       : IN    std_logic;
    SMA_MGT_TX_P     : OUT   std_logic;
    SMA_MGT_TX_N     : OUT   std_logic;
    SMA_MGT_RX_P     : IN    std_logic;
    SMA_MGT_RX_N     : IN    std_logic;
    --
    I2C_SCL          : INOUT std_logic;
    I2C_SDA          : INOUT std_logic;
    -- TE0741 B2B connector
    B12_L_P          : INOUT std_logic_vector(25 DOWNTO 0);
    B12_L_N          : INOUT std_logic_vector(25 DOWNTO 0);
    B13_L_P          : INOUT std_logic_vector(24 DOWNTO 0);
    B13_L_N          : INOUT std_logic_vector(24 DOWNTO 0);
    B14_L_P          : INOUT std_logic_vector(24 DOWNTO 0);
    B14_L_N          : INOUT std_logic_vector(24 DOWNTO 0);
    B15_L_P          : INOUT std_logic_vector(23 DOWNTO 0);
    B15_L_N          : INOUT std_logic_vector(23 DOWNTO 0);
    B16_L_P          : INOUT std_logic_vector(23 DOWNTO 0);
    B16_L_N          : INOUT std_logic_vector(23 DOWNTO 0)
  );
END top;

ARCHITECTURE Behavioral OF top IS
  -- Components
  COMPONENT global_clock_reset
    PORT (
      SYS_CLK_P  : IN  std_logic;
      SYS_CLK_N  : IN  std_logic;
      FORCE_RST  : IN  std_logic;
      -- output
      GLOBAL_RST : OUT std_logic;
      SYS_CLK    : OUT std_logic;
      LOCKED     : OUT std_logic;
      CLK_OUT1   : OUT std_logic;
      CLK_OUT2   : OUT std_logic;
      CLK_OUT3   : OUT std_logic;
      CLK_OUT4   : OUT std_logic
    );
  END COMPONENT;
  ---------------------------------------------< ten_gig_eth
  COMPONENT ten_gig_eth
    PORT (
      REFCLK_P             : IN  std_logic;  -- 156.25MHz for transceiver
      REFCLK_N             : IN  std_logic;
      RESET                : IN  std_logic;
      SFP_TX_P             : OUT std_logic;
      SFP_TX_N             : OUT std_logic;
      SFP_RX_P             : IN  std_logic;
      SFP_RX_N             : IN  std_logic;
      SFP_LOS              : IN  std_logic;  -- loss of receiver signal
      SFP_TX_DISABLE       : OUT std_logic;
      -- clk156.25 domain, clock generated by the core
      CLK156p25            : OUT std_logic;
      PCS_PMA_CORE_STATUS  : OUT std_logic_vector(7 DOWNTO 0);
      TX_STATISTICS_VECTOR : OUT std_logic_vector(25 DOWNTO 0);
      TX_STATISTICS_VALID  : OUT std_logic;
      RX_STATISTICS_VECTOR : OUT std_logic_vector(29 DOWNTO 0);
      RX_STATISTICS_VALID  : OUT std_logic;
      PAUSE_VAL            : IN  std_logic_vector(15 DOWNTO 0);
      PAUSE_REQ            : IN  std_logic;
      TX_IFG_DELAY         : IN  std_logic_vector(7 DOWNTO 0);
      -- emac control interface
      S_AXI_ACLK           : IN  std_logic;
      S_AXI_ARESETN        : IN  std_logic;
      S_AXI_AWADDR         : IN  std_logic_vector(10 DOWNTO 0);
      S_AXI_AWVALID        : IN  std_logic;
      S_AXI_AWREADY        : OUT std_logic;
      S_AXI_WDATA          : IN  std_logic_vector(31 DOWNTO 0);
      S_AXI_WVALID         : IN  std_logic;
      S_AXI_WREADY         : OUT std_logic;
      S_AXI_BRESP          : OUT std_logic_vector(1 DOWNTO 0);
      S_AXI_BVALID         : OUT std_logic;
      S_AXI_BREADY         : IN  std_logic;
      S_AXI_ARADDR         : IN  std_logic_vector(10 DOWNTO 0);
      S_AXI_ARVALID        : IN  std_logic;
      S_AXI_ARREADY        : OUT std_logic;
      S_AXI_RDATA          : OUT std_logic_vector(31 DOWNTO 0);
      S_AXI_RRESP          : OUT std_logic_vector(1 DOWNTO 0);
      S_AXI_RVALID         : OUT std_logic;
      S_AXI_RREADY         : IN  std_logic;
      -- tx_wr_clk domain
      TX_AXIS_FIFO_ARESETN : IN  std_logic;
      TX_AXIS_FIFO_ACLK    : IN  std_logic;
      TX_AXIS_FIFO_TDATA   : IN  std_logic_vector(63 DOWNTO 0);
      TX_AXIS_FIFO_TKEEP   : IN  std_logic_vector(7 DOWNTO 0);
      TX_AXIS_FIFO_TVALID  : IN  std_logic;
      TX_AXIS_FIFO_TLAST   : IN  std_logic;
      TX_AXIS_FIFO_TREADY  : OUT std_logic;
      -- rx_rd_clk domain
      RX_AXIS_FIFO_ARESETN : IN  std_logic;
      RX_AXIS_FIFO_ACLK    : IN  std_logic;
      RX_AXIS_FIFO_TDATA   : OUT std_logic_vector(63 DOWNTO 0);
      RX_AXIS_FIFO_TKEEP   : OUT std_logic_vector(7 DOWNTO 0);
      RX_AXIS_FIFO_TVALID  : OUT std_logic;
      RX_AXIS_FIFO_TLAST   : OUT std_logic;
      RX_AXIS_FIFO_TREADY  : IN  std_logic
    );
  END COMPONENT;
  COMPONENT ten_gig_eth_packet_gen
    PORT (
      RESET          : IN  std_logic;
      MEM_CLK        : IN  std_logic;
      MEM_WE         : IN  std_logic;   -- memory write enable
      MEM_ADDR       : IN  std_logic_vector(31 DOWNTO 0);
      MEM_D          : IN  std_logic_vector(31 DOWNTO 0);  -- memory data
      --
      TX_AXIS_ACLK   : IN  std_logic;
      TX_START       : IN  std_logic;
      TX_BYTES       : IN  std_logic_vector(15 DOWNTO 0);  -- number of bytes to send
      TX_AXIS_TDATA  : OUT std_logic_vector(63 DOWNTO 0);
      TX_AXIS_TKEEP  : OUT std_logic_vector(7 DOWNTO 0);
      TX_AXIS_TVALID : OUT std_logic;
      TX_AXIS_TLAST  : OUT std_logic;
      TX_AXIS_TREADY : IN  std_logic
    );
  END COMPONENT;
  COMPONENT ten_gig_eth_rx_parser
    PORT (
      RESET                : IN  std_logic;
      RX_AXIS_FIFO_ARESETN : OUT std_logic;
      -- Everything internal to this module is synchronous to this clock `ACLK'
      RX_AXIS_FIFO_ACLK    : IN  std_logic;
      RX_AXIS_FIFO_TDATA   : IN  std_logic_vector(63 DOWNTO 0);
      RX_AXIS_FIFO_TKEEP   : IN  std_logic_vector(7 DOWNTO 0);
      RX_AXIS_FIFO_TVALID  : IN  std_logic;
      RX_AXIS_FIFO_TLAST   : IN  std_logic;
      RX_AXIS_FIFO_TREADY  : OUT std_logic;
      -- Constants
      SRC_MAC              : IN  std_logic_vector(47 DOWNTO 0);
      SRC_IP               : IN  std_logic_vector(31 DOWNTO 0);
      SRC_PORT             : IN  std_logic_vector(15 DOWNTO 0);
      -- Command output fifo interface AFTER parsing the packet
      -- dstMAC(48) dstIP(32) dstPort(16) opcode(32)
      CMD_FIFO_Q           : OUT std_logic_vector(127 DOWNTO 0);
      CMD_FIFO_EMPTY       : OUT std_logic;
      CMD_FIFO_RDREQ       : IN  std_logic;
      CMD_FIFO_RDCLK       : IN  std_logic
    );
  END COMPONENT;
  ---------------------------------------------> ten_gig_eth
  ---------------------------------------------< gtx / aurora
  COMPONENT aurora_64b66b
    PORT (
      RESET               : IN  std_logic;
      SYS_CLK             : IN  std_logic;
      MGT_REFCLK_P        : IN  std_logic;
      MGT_REFCLK_N        : IN  std_logic;
      -- Data interfaces are synchronous to USER_CLK
      USER_CLK            : OUT std_logic;
      MGT_REFCLK_BUFG_OUT : OUT std_logic;
      -- TX AXI4 interface
      S_AXI_TX_TDATA      : IN  std_logic_vector(0 TO 63);
      S_AXI_TX_TVALID     : IN  std_logic;
      S_AXI_TX_TREADY     : OUT std_logic;
      -- RX AXI4 interface
      M_AXI_RX_TDATA      : OUT std_logic_vector(0 TO 63);
      M_AXI_RX_TVALID     : OUT std_logic;
      -- User flow control (UFC) TX
      UFC_TX_REQ          : IN  std_logic;
      S_AXI_UFC_TX_TDATA  : IN  std_logic_vector(0 TO 63);
      UFC_TX_MS           : IN  std_logic_vector(0 TO 7);
      S_AXI_UFC_TX_TVALID : IN  std_logic;
      S_AXI_UFC_TX_TREADY : OUT std_logic;
      -- UFC RX
      M_AXI_UFC_RX_TDATA  : OUT std_logic_vector(0 TO 63);
      M_AXI_UFC_RX_TKEEP  : OUT std_logic_vector(0 TO 7);
      M_AXI_UFC_RX_TLAST  : OUT std_logic;
      M_AXI_UFC_RX_TVALID : OUT std_logic;
      UFC_IN_PROGRESSn    : OUT std_logic;
      -- GTX pins
      RXP                 : IN  std_logic;
      RXN                 : IN  std_logic;
      TXP                 : OUT std_logic;
      TXN                 : OUT std_logic;
      -- Status
      STATUS              : OUT std_logic_vector(15 DOWNTO 0)
    );
  END COMPONENT;
  COMPONENT fifo_over_ufc
    GENERIC (
      FIFO_DATA_WIDTH   : positive := 32;
      AURORA_DATA_WIDTH : positive := 64
    );
    PORT (
      RESET            : IN  std_logic;
      AURORA_USER_CLK  : IN  std_logic;
      AURORA_TX_REQ    : OUT std_logic;
      AURORA_TX_MS     : OUT std_logic_vector(7 DOWNTO 0);
      AURORA_TX_TREADY : IN  std_logic;
      AURORA_TX_TDATA  : OUT std_logic_vector(AURORA_DATA_WIDTH-1 DOWNTO 0);
      AURORA_TX_TVALID : OUT std_logic;
      AURORA_RX_TDATA  : IN  std_logic_vector(AURORA_DATA_WIDTH-1 DOWNTO 0);
      AURORA_RX_TVALID : IN  std_logic;
      FIFO_CLK         : OUT std_logic;
      TX_FIFO_Q        : OUT std_logic_vector(FIFO_DATA_WIDTH-1 DOWNTO 0);
      TX_FIFO_WREN     : OUT std_logic;
      TX_FIFO_FULL     : IN  std_logic;
      RX_FIFO_Q        : IN  std_logic_vector(FIFO_DATA_WIDTH-1 DOWNTO 0);
      RX_FIFO_RDEN     : OUT std_logic;
      RX_FIFO_EMPTY    : IN  std_logic;
      ERR              : OUT std_logic
    );
  END COMPONENT;
  COMPONENT fifo36x512
    PORT (
      rst    : IN  std_logic;
      wr_clk : IN  std_logic;
      rd_clk : IN  std_logic;
      din    : IN  std_logic_vector(35 DOWNTO 0);
      wr_en  : IN  std_logic;
      rd_en  : IN  std_logic;
      dout   : OUT std_logic_vector(35 DOWNTO 0);
      full   : OUT std_logic;
      empty  : OUT std_logic
    );
  END COMPONENT;
  ---------------------------------------------> gtx / aurora
  ---------------------------------------------< UART/RS232
  COMPONENT control_interface
    PORT (
      RESET           : IN  std_logic;
      CLK             : IN  std_logic;    -- system clock
      -- From FPGA to PC
      FIFO_Q          : OUT std_logic_vector(35 DOWNTO 0);  -- interface fifo data output port
      FIFO_EMPTY      : OUT std_logic;    -- interface fifo "emtpy" signal
      FIFO_RDREQ      : IN  std_logic;    -- interface fifo read request
      FIFO_RDCLK      : IN  std_logic;    -- interface fifo read clock
      -- From PC to FPGA, FWFT
      CMD_FIFO_Q      : IN  std_logic_vector(35 DOWNTO 0);  -- interface command fifo data out port
      CMD_FIFO_EMPTY  : IN  std_logic;    -- interface command fifo "emtpy" signal
      CMD_FIFO_RDREQ  : OUT std_logic;    -- interface command fifo read request
      -- Digital I/O
      CONFIG_REG      : OUT std_logic_vector(511 DOWNTO 0); -- thirtytwo 16bit registers
      PULSE_REG       : OUT std_logic_vector(15 DOWNTO 0);  -- 16bit pulse register
      STATUS_REG      : IN  std_logic_vector(175 DOWNTO 0); -- eleven 16bit registers
      -- Memory interface
      MEM_WE          : OUT std_logic;    -- memory write enable
      MEM_ADDR        : OUT std_logic_vector(31 DOWNTO 0);
      MEM_DIN         : OUT std_logic_vector(31 DOWNTO 0);  -- memory data input
      MEM_DOUT        : IN  std_logic_vector(31 DOWNTO 0);  -- memory data output
      -- Data FIFO interface, FWFT
      DATA_FIFO_Q     : IN  std_logic_vector(31 DOWNTO 0);
      DATA_FIFO_EMPTY : IN  std_logic;
      DATA_FIFO_RDREQ : OUT std_logic;
      DATA_FIFO_RDCLK : OUT std_logic
    );
  END COMPONENT;
  ---------------------------------------------> UART/RS232
  ---------------------------------------------< I2C
  COMPONENT i2c_master
    GENERIC (
      INPUT_CLK_FREQENCY : integer := 100_000_000;
      -- BUS CLK freqency should be divided by multiples of 4 from input frequency
      BUS_CLK_FREQUENCY  : integer := 100_000
    );
    PORT (
      CLK       : IN  std_logic;        -- system clock 50Mhz
      RESET     : IN  std_logic;        -- active high reset
      START     : IN  std_logic;  -- rising edge triggers r/w; synchronous to CLK
      MODE      : IN  std_logic_vector(1 DOWNTO 0);  -- "00" : 1 bytes read or write, "01" : 2 bytes r/w, "10" : 3 bytes write only;
      SL_RW     : IN  std_logic;        -- '0' is write, '1' is read
      SL_ADDR   : IN  std_logic_vector(6 DOWNTO 0);  -- slave addr
      REG_ADDR  : IN  std_logic_vector(7 DOWNTO 0);  -- slave internal reg addr for read and write
      WR_DATA0  : IN  std_logic_vector(7 DOWNTO 0);  -- first data byte to write
      WR_DATA1  : IN  std_logic_vector(7 DOWNTO 0);  -- second data byte to write
      RD_DATA0  : OUT std_logic_vector(7 DOWNTO 0);  -- first data byte read
      RD_DATA1  : OUT std_logic_vector(7 DOWNTO 0);  -- second data byte read
      BUSY      : OUT std_logic;        -- indicates transaction in progress
      ACK_ERROR : OUT std_logic;        -- i2c has unexpected ack
      SDA_in    : IN  std_logic;        -- serial data input from i2c bus
      SDA_out   : OUT std_logic;        -- serial data output to i2c bus
      SDA_t     : OUT std_logic;  -- serial data direction to/from i2c bus, '1' is read-in
      SCL       : OUT std_logic         -- serial clock output to i2c bus
    );
  END COMPONENT;
  COMPONENT i2c_write_regmap
    GENERIC (
      REGMAP_FNAME        : string;
      INPUT_CLK_FREQENCY  : integer := 100_000_000;
      -- BUS CLK freqency should be divided by multiples of 4 from input frequency
      BUS_CLK_FREQUENCY   : integer := 100_000;
      START_DELAY_CYCLE   : integer := 100_000_000; -- ext_rst to happen # of clk cycles after START
      EXT_RST_WIDTH_CYCLE : integer := 1000;     -- pulse width of ext_rst in clk cycles
      EXT_RST_DELAY_CYCLE : integer := 100_000   -- 1st reg write to happen clk cycles after ext_rst
    );
    PORT (
      CLK       : IN  std_logic;        -- system clock 50Mhz
      RESET     : IN  std_logic;        -- active high reset
      START     : IN  std_logic;  -- rising edge triggers r/w; synchronous to CLK
      EXT_RSTn  : OUT std_logic;        -- active low for resetting the slave
      BUSY      : OUT std_logic;        -- indicates transaction in progress
      ACK_ERROR : OUT std_logic;        -- i2c has unexpected ack
      SDA_in    : IN  std_logic;        -- serial data input from i2c bus
      SDA_out   : OUT std_logic;        -- serial data output to i2c bus
      SDA_t     : OUT std_logic;  -- serial data direction to/from i2c bus, '1' is read-in
      SCL       : OUT std_logic         -- serial clock output to i2c bus
    );
  END COMPONENT;
  ---------------------------------------------> I2C
  ---------------------------------------------< shiftreg driver for DAC8568
  COMPONENT fifo2shiftreg
    GENERIC (
      DATA_WIDTH        : positive  := 32;  -- parallel data width
      CLK_DIV_WIDTH     : positive  := 16;
      DELAY_AFTER_SYNCn : natural   := 0;  -- number of SCLK cycles' wait after falling edge OF SYNCn
      SCLK_IDLE_LEVEL   : std_logic := '0';  -- High or Low for SCLK when not switching
      DOUT_DRIVE_EDGE   : std_logic := '1';  -- 1/0 rising/falling edge of SCLK drives new DOUT bit
      DIN_CAPTURE_EDGE  : std_logic := '0'  -- 1/0 rising/falling edge of SCLK captures new DIN bit
    );
    PORT (
      CLK      : IN  std_logic;         -- clock
      RESET    : IN  std_logic;         -- reset
      -- input data interface
      WR_CLK   : IN  std_logic;         -- FIFO write clock
      DINFIFO  : IN  std_logic_vector(15 DOWNTO 0);
      WR_EN    : IN  std_logic;
      WR_PULSE : IN  std_logic;  -- one pulse writes one word, regardless of pulse duration
      FULL     : OUT std_logic;
      -- captured data
      BUSY     : OUT std_logic;
      DATAOUT  : OUT std_logic_vector(DATA_WIDTH-1 DOWNTO 0);
      -- serial interface
      CLK_DIV  : IN  std_logic_vector(CLK_DIV_WIDTH-1 DOWNTO 0);  -- SCLK freq is CLK / 2**(CLK_DIV)
      SCLK     : OUT std_logic;
      DOUT     : OUT std_logic;
      SYNCn    : OUT std_logic;
      DIN      : IN  std_logic
    );
  END COMPONENT;
  ---------------------------------------------> shiftreg driver for DAC8568
  ---------------------------------------------< TMS serial io
  COMPONENT shiftreg_drive
    GENERIC (
      DATA_WIDTH        : positive  := 32;  -- parallel data width
      CLK_DIV_WIDTH     : positive  := 16;
      DELAY_AFTER_SYNCn : natural   := 0;  -- number of SCLK cycles' wait after falling edge OF SYNCn
      SCLK_IDLE_LEVEL   : std_logic := '0';  -- High or Low for SCLK when not switching
      DOUT_DRIVE_EDGE   : std_logic := '1';  -- 1/0 rising/falling edge of SCLK drives new DOUT bit
      DIN_CAPTURE_EDGE  : std_logic := '0'  -- 1/0 rising/falling edge of SCLK captures new DIN bit
    );
    PORT (
      CLK     : IN  std_logic;          -- clock
      RESET   : IN  std_logic;          -- reset
      -- internal data interface
      CLK_DIV : IN  std_logic_vector(CLK_DIV_WIDTH-1 DOWNTO 0);  -- SCLK freq is CLK / 2**(CLK_DIV)
      DATAIN  : IN  std_logic_vector(DATA_WIDTH-1 DOWNTO 0);
      START   : IN  std_logic;
      BUSY    : OUT std_logic;
      DATAOUT : OUT std_logic_vector(DATA_WIDTH-1 DOWNTO 0);
      -- external serial interface
      SCLK    : OUT std_logic;
      DOUT    : OUT std_logic;
      SYNCn   : OUT std_logic;
      DIN     : IN  std_logic
    );
  END COMPONENT;
  ---------------------------------------------> TMS serial io
  ---------------------------------------------< TMS SDM
  COMPONENT tms_sdm_recv
    GENERIC (
      NCH : positive := 19
    );
    PORT (
      RESET         : IN  std_logic;
      CLK           : IN  std_logic;  -- DELAY_* must be synchronous to this clock
      REFCLK        : IN  std_logic;    -- REFCLK (200MHz) for IDELAYCTRL
      DELAY_CHANNEL : IN  std_logic_vector(7 DOWNTO 0);  -- input iodelay channel selection
      DELAY_VALUE   : IN  std_logic_vector(4 DOWNTO 0);  -- input iodelay value
      DELAY_UPDATE  : IN  std_logic;    -- a pulse to update the delay value
      CLKFF_DIV     : IN  std_logic_vector(3 DOWNTO 0);
      CLKFF_P       : OUT std_logic;
      CLKFF_N       : OUT std_logic;
      CLK_LPBK_P    : IN  std_logic;
      CLK_LPBK_N    : IN  std_logic;
      CLK_LPBK      : OUT std_logic;
      SDM_OUT1_P    : IN  std_logic_vector(NCH-1 DOWNTO 0);
      SDM_OUT1_N    : IN  std_logic_vector(NCH-1 DOWNTO 0);
      SDM_OUT2_P    : IN  std_logic_vector(NCH-1 DOWNTO 0);
      SDM_OUT2_N    : IN  std_logic_vector(NCH-1 DOWNTO 0);
      DOUT          : OUT std_logic_vector(NCH*2-1 DOWNTO 0)
    );
  END COMPONENT;
  ---------------------------------------------> TMS SDM
  ---------------------------------------------< ADC, external, LTC2325-16
  COMPONENT adc_cnv_sipo
    GENERIC (
      NCH : positive := 20
    );
    PORT (
      RESET         : IN  std_logic;
      CLK           : IN  std_logic;  -- DELAY_* must be synchronous to this clock
      REFCLK        : IN  std_logic;    -- REFCLK (200MHz) for IDELAYCTRL
      DELAY_CHANNEL : IN  std_logic_vector(7 DOWNTO 0);  -- ADC data input iodelay channel selection
      DELAY_VALUE   : IN  std_logic_vector(4 DOWNTO 0);  -- ADC data input iodelay value
      DELAY_UPDATE  : IN  std_logic;    -- a pulse to update the delay value
      CLKFF_DIV     : IN  std_logic_vector(3 DOWNTO 0);
      CLKFF_P       : OUT std_logic;
      CLKFF_N       : OUT std_logic;
      CLK_LPBK_P    : IN  std_logic;
      CLK_LPBK_N    : IN  std_logic;
      CLK_LPBK      : OUT std_logic;
      CNV_N_P       : OUT std_logic;
      CNV_N_N       : OUT std_logic;
      CNV_N         : OUT std_logic;
      INPUTS_P      : IN  std_logic_vector(NCH-1 DOWNTO 0);
      INPUTS_N      : IN  std_logic_vector(NCH-1 DOWNTO 0);
      INPUTS_OUT    : OUT std_logic_vector(NCH-1 DOWNTO 0);
      DOUT          : OUT std_logic_vector(NCH*16-1 DOWNTO 0);
      DOUT_VALID    : OUT std_logic
    );
  END COMPONENT;
  ---------------------------------------------> ADC, external, LTC2325-16
  ---------------------------------------------< debug : ILA and VIO (`Chipscope')
  COMPONENT dbg_ila
    PORT (
      CLK    : IN std_logic;
      PROBE0 : IN std_logic_vector(63 DOWNTO 0);
      PROBE1 : IN std_logic_vector(79 DOWNTO 0);
      PROBE2 : IN std_logic_vector(79 DOWNTO 0);
      PROBE3 : IN std_logic_vector(2047 DOWNTO 0)
    );
  END COMPONENT;
  COMPONENT dbg_ila1
    PORT (
      CLK    : IN std_logic;
      PROBE0 : IN std_logic_vector(15 DOWNTO 0);
      PROBE1 : IN std_logic_vector(15 DOWNTO 0)
    );
  END COMPONENT;
  COMPONENT dbg_vio
    PORT (
      CLK        : IN  std_logic;
      PROBE_IN0  : IN  std_logic_vector(63 DOWNTO 0);
      PROBE_IN1  : IN  std_logic_vector(63 DOWNTO 0);
      PROBE_IN2  : IN  std_logic_vector(63 DOWNTO 0);
      PROBE_IN3  : IN  std_logic_vector(63 DOWNTO 0);
      PROBE_IN4  : IN  std_logic_vector(63 DOWNTO 0);
      PROBE_IN5  : IN  std_logic_vector(63 DOWNTO 0);
      PROBE_IN6  : IN  std_logic_vector(63 DOWNTO 0);
      PROBE_IN7  : IN  std_logic_vector(63 DOWNTO 0);
      PROBE_IN8  : IN  std_logic_vector(35 DOWNTO 0);
      PROBE_OUT0 : OUT std_logic_vector(63 DOWNTO 0)
    );
  END COMPONENT;
  ---------------------------------------------> debug : ILA and VIO (`Chipscope')

  -- Signals
  SIGNAL reset                             : std_logic;
  SIGNAL sys_clk                           : std_logic;
  SIGNAL global_clk_locked                 : std_logic;
  SIGNAL clk_50MHz                         : std_logic;
  SIGNAL clk_100MHz                        : std_logic;
  SIGNAL clk_125MHz                        : std_logic;
  SIGNAL clk_200MHz                        : std_logic;
  SIGNAL clk_250MHz                        : std_logic;
  SIGNAL clk_sgmii_i                       : std_logic;
  SIGNAL clk_sgmii                         : std_logic;
  SIGNAL clk156p25                         : std_logic;
  SIGNAL clk_user                          : std_logic;
  ---------------------------------------------< UART/RS232
  SIGNAL uart_rx_data                      : std_logic_vector(7 DOWNTO 0);
  SIGNAL uart_rx_rdy                       : std_logic;
  SIGNAL control_clk                       : std_logic;
  SIGNAL control_fifo_q                    : std_logic_vector(35 DOWNTO 0);
  SIGNAL control_fifo_rdreq                : std_logic;
  SIGNAL control_fifo_empty                : std_logic;
  SIGNAL control_fifo_rdclk                : std_logic;
  SIGNAL cmd_fifo_q                        : std_logic_vector(35 DOWNTO 0);
  SIGNAL cmd_fifo_empty                    : std_logic;
  SIGNAL cmd_fifo_rdreq                    : std_logic;
  -- thirtytwo 16bit registers
  SIGNAL config_reg                        : std_logic_vector(511 DOWNTO 0);
  -- 16bit pulse register
  SIGNAL pulse_reg                         : std_logic_vector(15 DOWNTO 0);
  -- eleven 16bit registers
  SIGNAL status_reg                        : std_logic_vector(175 DOWNTO 0) := (OTHERS => '0');
  SIGNAL control_mem_we                    : std_logic;
  SIGNAL control_mem_addr                  : std_logic_vector(31 DOWNTO 0);
  SIGNAL control_mem_din                   : std_logic_vector(31 DOWNTO 0);
  ---------------------------------------------> UART/RS232
  ---------------------------------------------< gtx / aurora
  SIGNAL aurora_reset                      : std_logic;
  SIGNAL aurora_status                     : std_logic_vector(15 DOWNTO 0);
  SIGNAL aurora_user_clk                   : std_logic;
  SIGNAL aurora_ufc_tx_req                 : std_logic;
  SIGNAL aurora_ufc_tx_tdata               : std_logic_vector(63 DOWNTO 0);
  SIGNAL aurora_ufc_tx_ms                  : std_logic_vector(7 DOWNTO 0);
  SIGNAL aurora_ufc_tx_tvalid              : std_logic;
  SIGNAL aurora_ufc_tx_tready              : std_logic;
  SIGNAL aurora_ufc_rx_tdata               : std_logic_vector(63 DOWNTO 0);
  SIGNAL aurora_ufc_rx_tkeep               : std_logic_vector(7 DOWNTO 0);
  SIGNAL aurora_ufc_rx_tlast               : std_logic;
  SIGNAL aurora_ufc_rx_tvalid              : std_logic;
  SIGNAL aurora_ufc_in_progress_n          : std_logic;
  SIGNAL aurora_ufc_tx_fifo_q              : std_logic_vector(31 DOWNTO 0);
  SIGNAL aurora_ufc_tx_fifo_wren           : std_logic;
  SIGNAL aurora_ufc_tx_fifo_full           : std_logic;
  SIGNAL aurora_tx_tdata                   : std_logic_vector(63 DOWNTO 0);
  SIGNAL aurora_tx_tvalid                  : std_logic;
  SIGNAL aurora_tx_tready                  : std_logic;
  SIGNAL aurora_rx_tdata                   : std_logic_vector(63 DOWNTO 0);
  SIGNAL aurora_rx_tvalid                  : std_logic;
  ---------------------------------------------> gtx / aurora
  ---------------------------------------------< ten_gig_eth
  SIGNAL sfp_tx_disable_i                  : std_logic;
  SIGNAL sPcs_pma_core_status              : std_logic_vector(7 DOWNTO 0);
  SIGNAL sEmac_status_vector               : std_logic_vector(1 DOWNTO 0);
  SIGNAL sTx_axis_fifo_aresetn             : std_logic;
  SIGNAL sTx_axis_fifo_aclk                : std_logic;
  SIGNAL sTx_axis_fifo_tdata               : std_logic_vector(63 DOWNTO 0);
  SIGNAL sTx_axis_fifo_tkeep               : std_logic_vector(7 DOWNTO 0);
  SIGNAL sTx_axis_fifo_tvalid              : std_logic;
  SIGNAL sTx_axis_fifo_tlast               : std_logic;
  SIGNAL sTx_axis_fifo_tready              : std_logic;
  SIGNAL sRx_axis_fifo_aresetn             : std_logic;
  SIGNAL sRx_axis_fifo_aclk                : std_logic;
  SIGNAL sRx_axis_fifo_tdata               : std_logic_vector(63 DOWNTO 0);
  SIGNAL sRx_axis_fifo_tkeep               : std_logic_vector(7 DOWNTO 0);
  SIGNAL sRx_axis_fifo_tvalid              : std_logic;
  SIGNAL sRx_axis_fifo_tlast               : std_logic;
  SIGNAL sRx_axis_fifo_tready              : std_logic;
  -- control interface
  SIGNAL s_axi_aclk                        : std_logic;
  SIGNAL s_axi_aresetn                     : std_logic;
  SIGNAL s_axi_awaddr                      : std_logic_vector(10 DOWNTO 0);
  SIGNAL s_axi_awvalid                     : std_logic;
  SIGNAL s_axi_awready                     : std_logic;
  SIGNAL s_axi_wdata                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL s_axi_wvalid                      : std_logic;
  SIGNAL s_axi_wready                      : std_logic;
  SIGNAL s_axi_bresp                       : std_logic_vector(1 DOWNTO 0);
  SIGNAL s_axi_bvalid                      : std_logic;
  SIGNAL s_axi_bready                      : std_logic;
  SIGNAL s_axi_araddr                      : std_logic_vector(10 DOWNTO 0);
  SIGNAL s_axi_arvalid                     : std_logic;
  SIGNAL s_axi_arready                     : std_logic;
  SIGNAL s_axi_rdata                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL s_axi_rresp                       : std_logic_vector(1 DOWNTO 0);
  SIGNAL s_axi_rvalid                      : std_logic;
  SIGNAL s_axi_rready                      : std_logic;
  -- packets
  SIGNAL ten_gig_eth_tx_start              : std_logic;
  SIGNAL tge_cmd_fifo_q                    : std_logic_vector(127 DOWNTO 0);
  SIGNAL tge_cmd_fifo_empty                : std_logic;
  SIGNAL tge_cmd_fifo_rdreq                : std_logic;
  ---------------------------------------------> ten_gig_eth
  SIGNAL usr_data_output                   : std_logic_vector (7 DOWNTO 0);
  ---------------------------------------------< IDATA
  SIGNAL TRIG_OUT_0                        : std_logic;
  SIGNAL idata_cmd_out                     : std_logic_vector(63 DOWNTO 0);
  SIGNAL idata_cmd_out_val                 : std_logic;
  SIGNAL idata_cmd_in                      : std_logic_vector(63 DOWNTO 0);
  SIGNAL idata_cmd_in_val                  : std_logic;
  SIGNAL idata_adc_data_clk                : std_logic;
  SIGNAL idata_adc_refout_clkdiv           : std_logic;
  SIGNAL idata_adc_data0                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data1                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data2                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data3                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data4                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data5                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data6                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data7                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data8                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data9                   : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data10                  : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_adc_data11                  : std_logic_vector(15 DOWNTO 0);
  SIGNAL idata_data_fifo_reset             : std_logic;
  SIGNAL idata_data_fifo_rdclk             : std_logic;
  SIGNAL idata_data_fifo_din               : std_logic_vector(255 DOWNTO 0);
  SIGNAL idata_channel_avg_outdata_q       : std_logic_vector(255 DOWNTO 0);
  SIGNAL idata_channel_avg_outvalid        : std_logic;
  SIGNAL idata_data_fifo_wren              : std_logic;
  SIGNAL idata_data_fifo_rden              : std_logic;
  SIGNAL idata_data_fifo_dout              : std_logic_vector(31 DOWNTO 0);
  SIGNAL idata_data_fifo_full              : std_logic;
  SIGNAL idata_data_fifo_empty             : std_logic;
  SIGNAL idata_idata_fifo_q                : std_logic_vector(255 DOWNTO 0);
  SIGNAL idata_idata_fifo_wren             : std_logic;
  SIGNAL idata_idata_fifo_rden             : std_logic;
  SIGNAL idata_idata_fifo_full             : std_logic;
  SIGNAL idata_idata_fifo_empty            : std_logic;
  SIGNAL idata_trig_allow                  : std_logic;
  SIGNAL idata_trig_in                     : std_logic;
  SIGNAL idata_trig_synced                 : std_logic;
  SIGNAL idata_data_wr_start               : std_logic;
  SIGNAL idata_data_wr_busy                : std_logic;
  SIGNAL idata_data_wr_wrapped             : std_logic;
  ---------------------------------------------> IDATA
  ---------------------------------------------< I2C
  SIGNAL i2c_sda_out                       : std_logic;
  SIGNAL i2c_sda_in                        : std_logic;
  SIGNAL i2c_sda_t                         : std_logic;
  SIGNAL i2c_scl_out                       : std_logic;
  SIGNAL i2c1_sda_out                      : std_logic;
  SIGNAL i2c1_sda_in                       : std_logic;
  SIGNAL i2c1_sda_t                        : std_logic;
  SIGNAL i2c1_scl_out                      : std_logic;
  ---------------------------------------------> I2C
  ---------------------------------------------< shiftreg driver for DAC8568
  SIGNAL spi_sclk                          : std_logic;
  SIGNAL spi_dout                          : std_logic;
  SIGNAL spi_sync_n                        : std_logic;
  SIGNAL spi_din                           : std_logic;
  ---------------------------------------------> shiftreg driver for DAC8568
  ---------------------------------------------< TMS
  SIGNAL tms_pwr_on                        : std_logic;
  SIGNAL tms_sio_a                         : std_logic_vector(2 DOWNTO 0);
  SIGNAL tms_sdi                           : std_logic;
  SIGNAL tms_sdo                           : std_logic;
  SIGNAL tms_sck                           : std_logic;
  SIGNAL dac_din                           : std_logic;
  SIGNAL dac_sclk                          : std_logic;
  SIGNAL dac_sync_n                        : std_logic;
  SIGNAL tms_reset                         : std_logic;
  SIGNAL tms_sdm_clk_src_sel               : std_logic;
  SIGNAL tms_sdm_clkff_div                 : std_logic_vector(3 DOWNTO 0);
  SIGNAL tms_sdm_clk_lpbk                  : std_logic;
  SIGNAL tms_sdm_out1_p                    : std_logic_vector(18 DOWNTO 0);
  SIGNAL tms_sdm_out1_n                    : std_logic_vector(18 DOWNTO 0);
  SIGNAL tms_sdm_out2_p                    : std_logic_vector(18 DOWNTO 0);
  SIGNAL tms_sdm_out2_n                    : std_logic_vector(18 DOWNTO 0);
  SIGNAL tms_sdm_out                       : std_logic_vector(37 DOWNTO 0);
  SIGNAL adc_clk_src_sel                   : std_logic;
  SIGNAL adc_clkff_div                     : std_logic_vector(3 DOWNTO 0);
  SIGNAL adc_clk0_lpbk                     : std_logic;
  SIGNAL adc_sdrn_ddr                      : std_logic;
  SIGNAL adc_cnv_n                         : std_logic;
  SIGNAL adc_sdo_p                         : std_logic_vector(19 DOWNTO 0);
  SIGNAL adc_sdo_n                         : std_logic_vector(19 DOWNTO 0);
  SIGNAL adc_sdo                           : std_logic_vector(19 DOWNTO 0);
  SIGNAL adc_dout                          : std_logic_vector(20*16-1 DOWNTO 0);
  SIGNAL adc_dout_valid                    : std_logic;
  ---------------------------------------------> TMS
  ---------------------------------------------< debug
  SIGNAL dbg_ila_probe0                           : std_logic_vector(63 DOWNTO 0);
  SIGNAL dbg_ila_probe1                           : std_logic_vector(79 DOWNTO 0);
  SIGNAL dbg_ila_probe2                           : std_logic_vector(79 DOWNTO 0);
  SIGNAL dbg_ila_probe3                           : std_logic_vector(2047 DOWNTO 0);
  SIGNAL dbg_vio_probe_out0                       : std_logic_vector(63 DOWNTO 0);
  SIGNAL dbg_ila1_probe0                          : std_logic_vector(15 DOWNTO 0);
  SIGNAL dbg_ila1_probe1                          : std_logic_vector(15 DOWNTO 0);
  ATTRIBUTE mark_debug                            : string;
  ATTRIBUTE keep                                  : string;
  ATTRIBUTE mark_debug OF uart_rx_data            : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF uart_rx_rdy             : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF cmd_fifo_q              : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF cmd_fifo_empty          : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF cmd_fifo_rdreq          : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF config_reg              : SIGNAL IS "true";
--ATTRIBUTE mark_debug OF status_reg              : SIGNAL IS "true";
--ATTRIBUTE mark_debug OF pulse_reg               : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF control_mem_we          : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF control_mem_addr        : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF control_mem_din         : SIGNAL IS "true";
  --
  ATTRIBUTE mark_debug OF sPcs_pma_core_status    : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sEmac_status_vector     : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sTx_axis_fifo_aresetn   : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sTx_axis_fifo_aclk      : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sTx_axis_fifo_tdata     : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sTx_axis_fifo_tkeep     : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sTx_axis_fifo_tvalid    : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sTx_axis_fifo_tlast     : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sTx_axis_fifo_tready    : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sRx_axis_fifo_aresetn   : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sRx_axis_fifo_aclk      : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sRx_axis_fifo_tdata     : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sRx_axis_fifo_tkeep     : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sRx_axis_fifo_tvalid    : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sRx_axis_fifo_tlast     : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF sRx_axis_fifo_tready    : SIGNAL IS "true";
  --ATTRIBUTE mark_debug OF ten_gig_eth_tx_start    : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF tge_cmd_fifo_q          : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF tge_cmd_fifo_empty      : SIGNAL IS "true";
  ATTRIBUTE mark_debug OF tge_cmd_fifo_rdreq      : SIGNAL IS "true";
  ---------------------------------------------> debug

BEGIN
  ---------------------------------------------< Clock
  global_clock_reset_inst : global_clock_reset
    PORT MAP (
      SYS_CLK_P  => SYS_CLK_P,
      SYS_CLK_N  => SYS_CLK_N,
      FORCE_RST  => SYS_RST,
      -- output
      GLOBAL_RST => reset,
      SYS_CLK    => sys_clk,
      LOCKED     => global_clk_locked,
      CLK_OUT1   => clk_50MHz,
      CLK_OUT2   => OPEN,
      CLK_OUT3   => OPEN,
      CLK_OUT4   => clk_200MHz
    );
  clk_100MHz <= sys_clk;

  -- user_clk_ibufds_inst : IBUFDS
  --   GENERIC MAP (
  --     DIFF_TERM    => true,             -- Differential Termination
  --     IBUF_LOW_PWR => false,  -- Low power (TRUE) vs. performance (FALSE) setting for referenced I/O standards
  --     IOSTANDARD   => "LVDS"
  --   )
  --   PORT MAP (
  --     O  => clk_user,                   -- Buffer output
  --     I  => USER_CLK_P,  -- Diff_p buffer input (connect directly to top-level port)
  --     IB => USER_CLK_N   -- Diff_n buffer input (connect directly to top-level port)
  --   );

  -- gtx/gth reference clock can be used as general purpose clock this way
  -- sgmiiclk_ibufds_inst : IBUFDS_GTE2
  --   PORT MAP (
  --     O     => clk_sgmii_i,
  --     ODIV2 => OPEN,
  --     CEB   => '0',
  --     I     => SGMIICLK_Q0_P,
  --     IB    => SGMIICLK_Q0_N
  --   );
  -- sgmiiclk_bufg_inst : BUFG
  --   PORT MAP (
  --     I => clk_sgmii_i,
  --     O => clk_sgmii
  --   );
  clk_125MHz <= clk_sgmii;
  ---------------------------------------------> Clock
  ---------------------------------------------< debug : ILA and VIO (`Chipscope')
  dbg_cores : IF ENABLE_DEBUG GENERATE
    dbg_ila_inst : dbg_ila
      PORT MAP (
        CLK    => sys_clk,
        PROBE0 => dbg_ila_probe0,
        PROBE1 => dbg_ila_probe1,
        PROBE2 => dbg_ila_probe2,
        PROBE3 => dbg_ila_probe3
      );
    dbg_vio_inst : dbg_vio
      PORT MAP (
        CLK        => sys_clk,
        PROBE_IN0  => config_reg(64*1-1 DOWNTO 64*0),
        PROBE_IN1  => config_reg(64*2-1 DOWNTO 64*1),
        PROBE_IN2  => config_reg(64*3-1 DOWNTO 64*2),
        PROBE_IN3  => config_reg(64*4-1 DOWNTO 64*3),
        PROBE_IN4  => config_reg(64*5-1 DOWNTO 64*4),
        PROBE_IN5  => config_reg(64*6-1 DOWNTO 64*5),
        PROBE_IN6  => config_reg(64*7-1 DOWNTO 64*6),
        PROBE_IN7  => x"00000000000000" & sPcs_pma_core_status, -- config_reg(64*8-1 DOWNTO 64*7),
        PROBE_IN8  => cmd_fifo_q,
        PROBE_OUT0 => dbg_vio_probe_out0
      );
    --dbg_ila1_inst : dbg_ila1
    --  PORT MAP (
    --    CLK    => sys_clk,
    --    PROBE0 => dbg_ila1_probe0,
    --    PROBE1 => dbg_ila1_probe1
    --  );
  END GENERATE dbg_cores;
  ---------------------------------------------> debug : ILA and VIO (`Chipscope')
  ---------------------------------------------< UART/RS232
  uart_cores : IF false GENERATE
    uartio_inst : uartio
      GENERIC MAP (
        -- tick repetition frequency is (input freq) / (2**COUNTER_WIDTH / DIVISOR)
        COUNTER_WIDTH => 16,
        DIVISOR       => 1208*2
      )
      PORT MAP (
        CLK     => clk_50MHz,
        RESET   => reset,
        RX_DATA => uart_rx_data,
        RX_RDY  => uart_rx_rdy,
        TX_DATA => x"00",
        TX_EN   => '1',
        TX_RDY  => dbg_ila_probe0(2),
        -- serial lines
        RX_PIN  => '0',
        TX_PIN  => OPEN
      );

    --dbg_ila1_probe0(7 DOWNTO 0)  <= uart_rx_data;
    --dbg_ila1_probe0(8)           <= uart_rx_rdy;
    --dbg_ila1_probe0(9)           <= USB_TX;

    -- dbg_ila_probe0(63 DOWNTO 32) <= cmd_fifo_q(31 DOWNTO 0);
    dbg_ila_probe0(31)           <= cmd_fifo_empty;
    dbg_ila_probe0(30)           <= cmd_fifo_rdreq;

    byte2cmd_inst : byte2cmd
      PORT MAP (
        CLK            => clk_50MHz,
        RESET          => reset,
        -- byte in
        RX_DATA        => uart_rx_data,
        RX_RDY         => uart_rx_rdy,
        -- cmd out
        CMD_FIFO_Q     => OPEN,-- cmd_fifo_q,
        CMD_FIFO_EMPTY => OPEN,-- cmd_fifo_empty,
        CMD_FIFO_RDCLK => control_clk,
        CMD_FIFO_RDREQ => '0'  -- cmd_fifo_rdreq
      );
  END GENERATE uart_cores;

  control_clk <= clk_100MHz;
  control_interface_inst : control_interface
    PORT MAP (
      RESET => reset,
      CLK   => control_clk,
      -- From FPGA to PC
      FIFO_Q          => control_fifo_q,
      FIFO_EMPTY      => control_fifo_empty,
      FIFO_RDREQ      => control_fifo_rdreq,
      FIFO_RDCLK      => control_fifo_rdclk,
      -- From PC to FPGA, FWFT
      CMD_FIFO_Q      => cmd_fifo_q,
      CMD_FIFO_EMPTY  => cmd_fifo_empty,
      CMD_FIFO_RDREQ  => cmd_fifo_rdreq,
      -- Digital I/O
      CONFIG_REG      => config_reg,
      PULSE_REG       => pulse_reg,
      STATUS_REG      => status_reg,
      -- Memory interface
      MEM_WE          => control_mem_we,
      MEM_ADDR        => control_mem_addr,
      MEM_DIN         => control_mem_din,
      MEM_DOUT        => (OTHERS => '0'),
      -- Data FIFO interface, FWFT
      DATA_FIFO_Q     => idata_data_fifo_dout,
      DATA_FIFO_EMPTY => idata_data_fifo_empty,
      DATA_FIFO_RDREQ => idata_data_fifo_rden,
      DATA_FIFO_RDCLK => idata_data_fifo_rdclk
    );
  dbg_ila_probe0(18 DOWNTO 3) <= pulse_reg;
  ---------------------------------------------> UART/RS232
  ---------------------------------------------< ten_gig_eth
  B14_L_N(5)  <= '1';                   -- TE0741 CLK_EN
  B14_L_N(21) <= '1';                   -- TE0741 EN_MGT
  ten_gig_eth_cores : IF ENABLE_TEN_GIG_ETH GENERATE
    ten_gig_eth_inst : ten_gig_eth
      PORT MAP (
        REFCLK_P             => MGT_CLK3_P, -- 156.25MHz for transceiver
        REFCLK_N             => MGT_CLK3_N,
        RESET                => reset,
        SFP_TX_P             => SFP_TX_P,
        SFP_TX_N             => SFP_TX_N,
        SFP_RX_P             => SFP_RX_P,
        SFP_RX_N             => SFP_RX_N,
        SFP_LOS              => SFP_LOS_LS,  -- loss of receiver signal
        SFP_TX_DISABLE       => sfp_tx_disable_i,
        -- clk156.25 domain, clock generated by the core
        CLK156p25            => clk156p25,
        PCS_PMA_CORE_STATUS  => sPcs_pma_core_status,
        TX_STATISTICS_VECTOR => OPEN,
        TX_STATISTICS_VALID  => OPEN,
        RX_STATISTICS_VECTOR => OPEN,
        RX_STATISTICS_VALID  => OPEN,
        PAUSE_VAL            => (OTHERS => '0'),
        PAUSE_REQ            => '0',
        TX_IFG_DELAY         => x"ff",
        -- emac control interface
        S_AXI_ACLK           => s_axi_aclk,
        S_AXI_ARESETN        => s_axi_aresetn,
        S_AXI_AWADDR         => s_axi_awaddr,
        S_AXI_AWVALID        => s_axi_awvalid,
        S_AXI_AWREADY        => s_axi_awready,
        S_AXI_WDATA          => s_axi_wdata,
        S_AXI_WVALID         => s_axi_wvalid,
        S_AXI_WREADY         => s_axi_wready,
        S_AXI_BRESP          => s_axi_bresp,
        S_AXI_BVALID         => s_axi_bvalid,
        S_AXI_BREADY         => s_axi_bready,
        S_AXI_ARADDR         => s_axi_araddr,
        S_AXI_ARVALID        => s_axi_arvalid,
        S_AXI_ARREADY        => s_axi_arready,
        S_AXI_RDATA          => s_axi_rdata,
        S_AXI_RRESP          => s_axi_rresp,
        S_AXI_RVALID         => s_axi_rvalid,
        S_AXI_RREADY         => s_axi_rready,
        -- tx_wr_clk domain
        TX_AXIS_FIFO_ARESETN => sTx_axis_fifo_aresetn,
        Tx_AXIS_FIFO_ACLK    => sTx_axis_fifo_aclk,
        TX_AXIS_FIFO_TDATA   => sTx_axis_fifo_tdata,
        TX_AXIS_FIFO_TKEEP   => sTx_axis_fifo_tkeep,
        TX_AXIS_FIFO_TVALID  => sTx_axis_fifo_tvalid,
        TX_AXIS_FIFO_TLAST   => sTx_axis_fifo_tlast,
        TX_AXIS_FIFO_TREADY  => sTx_axis_fifo_tready,
        -- rx_rd_clk domain
        RX_AXIS_FIFO_ARESETN => sRx_axis_fifo_aresetn,
        RX_AXIS_FIFO_ACLK    => sRx_axis_fifo_aclk,
        RX_AXIS_FIFO_TDATA   => sRx_axis_fifo_tdata,
        RX_AXIS_FIFO_TKEEP   => sRx_axis_fifo_tkeep,
        RX_AXIS_FIFO_TVALID  => sRx_axis_fifo_tvalid,
        RX_AXIS_FIFO_TLAST   => sRx_axis_fifo_tlast,
        RX_AXIS_FIFO_TREADY  => sRx_axis_fifo_tready
      );

    SFP_TX_DISABLE_N   <= NOT sfp_tx_disable_i;
    LED8Bit(7)         <= sPcs_pma_core_status(0);
    LED8Bit(6)         <= NOT sfp_tx_disable_i;
    LED8Bit(5)         <= NOT SFP_LOS_LS;
    s_axi_aclk         <= clk_50MHz;
    sTx_axis_fifo_aclk <= clk_200MHz;
    sRx_axis_fifo_aclk <= sTx_axis_fifo_aclk;

    s_axi_aresetn         <= '1';
    sTx_axis_fifo_aresetn <= '1';
    -- sRx_axis_fifo_aresetn <= '1';

    ten_gig_eth_packet_gen_inst : ten_gig_eth_packet_gen
      PORT MAP (
        RESET          => reset,
        MEM_CLK        => control_clk,
        MEM_WE         => control_mem_we,
        MEM_ADDR       => control_mem_addr,
        MEM_D          => control_mem_din,
        --
        TX_AXIS_ACLK   => sTx_axis_fifo_aclk,
        TX_START       => ten_gig_eth_tx_start,
        TX_BYTES       => config_reg(15 DOWNTO 0),
        TX_AXIS_TDATA  => OPEN, -- sTx_axis_fifo_tdata,
        TX_AXIS_TKEEP  => sTx_axis_fifo_tkeep,
        TX_AXIS_TVALID => sTx_axis_fifo_tvalid,
        TX_AXIS_TLAST  => sTx_axis_fifo_tlast,
        TX_AXIS_TREADY => sTx_axis_fifo_tready
      );

    ten_gig_eth_rx_parser_inst : ten_gig_eth_rx_parser
      PORT MAP (
        RESET                => reset,
        RX_AXIS_FIFO_ARESETN => sRx_axis_fifo_aresetn,
        -- Everything internal to this module is synchronous to this clock `ACLK'
        RX_AXIS_FIFO_ACLK    => sRx_axis_fifo_aclk,
        RX_AXIS_FIFO_TDATA   => sRx_axis_fifo_tdata,
        RX_AXIS_FIFO_TKEEP   => sRx_axis_fifo_tkeep,
        RX_AXIS_FIFO_TVALID  => sRx_axis_fifo_tvalid,
        RX_AXIS_FIFO_TLAST   => sRx_axis_fifo_tlast,
        RX_AXIS_FIFO_TREADY  => sRx_axis_fifo_tready,
        -- Constants
        SRC_MAC              => x"000a3502a759",
        SRC_IP               => x"c0a80302",
        SRC_PORT             => x"ea62",
        -- Command output fifo interface AFTER parsing the packet
        -- dstMAC(48) dstIP(32) dstPort(16) opcode(32)
        CMD_FIFO_Q           => tge_cmd_fifo_q,
        CMD_FIFO_EMPTY       => tge_cmd_fifo_empty,
        CMD_FIFO_RDREQ       => '1',
        CMD_FIFO_RDCLK       => clk_200MHz
      );

    ten_gig_eth_tx_start <= pulse_reg(0);

    dbg_ila_probe0(0) <= clk156p25;
    dbg_ila_probe0(1) <= ten_gig_eth_tx_start;

    dbg_ila_probe1(79 DOWNTO 16) <= sTx_axis_fifo_tdata;
    dbg_ila_probe1(15 DOWNTO 8)  <= sTx_axis_fifo_tkeep;
    dbg_ila_probe1(7)            <= sTx_axis_fifo_tvalid;
    dbg_ila_probe1(6)            <= sTx_axis_fifo_tlast;
    dbg_ila_probe1(5)            <= sTx_axis_fifo_tready;
    --dbg_ila_probe2(79 DOWNTO 16) <= sRx_axis_fifo_tdata;
    --dbg_ila_probe2(79 DOWNTO 48) <= control_mem_addr;
    --dbg_ila_probe2(47 DOWNTO 16) <= control_mem_din;
    --dbg_ila_probe2(15 DOWNTO 8)  <= sRx_axis_fifo_tkeep;
    dbg_ila_probe2(7)            <= sRx_axis_fifo_tvalid;
    dbg_ila_probe2(6)            <= sRx_axis_fifo_tlast;
    dbg_ila_probe2(5)            <= sRx_axis_fifo_tready;
    dbg_ila_probe2(4)            <= control_mem_we;
    --
    --dbg_ila_probe3(127 DOWNTO 0) <= tge_cmd_fifo_q;
    --dbg_ila_probe3(128)          <= tge_cmd_fifo_empty;
  END GENERATE ten_gig_eth_cores;
  ---------------------------------------------> ten_gig_eth
  ---------------------------------------------< gtx / aurora
  -- SFP_TX_DISABLE_N <= '1';
  -- LED8Bit(0) <= NOT B14_L_P(19);        -- NOT SFP_LOS_LS;  -- SFP is plugged in.
  LED8Bit(1) <= aurora_status(0);                           -- link up
  aurora_64b66b_inst : aurora_64b66b
    PORT MAP (
      RESET               => aurora_reset,
      SYS_CLK             => clk_100MHz,
      MGT_REFCLK_P        => SGMIICLK_Q0_P,
      MGT_REFCLK_N        => SGMIICLK_Q0_N,
      -- Data interfaces are synchronous to USER_CLK
      USER_CLK            => aurora_user_clk,
      MGT_REFCLK_BUFG_OUT => clk_sgmii,
      -- TX AXI4 interface
      S_AXI_TX_TDATA      => aurora_tx_tdata,
      S_AXI_TX_TVALID     => aurora_tx_tvalid,
      S_AXI_TX_TREADY     => aurora_tx_tready,
      -- RX AXI4 interface
      M_AXI_RX_TDATA      => aurora_rx_tdata,
      M_AXI_RX_TVALID     => aurora_rx_tvalid,
      -- User flow control (UFC) TX
      UFC_TX_REQ          => aurora_ufc_tx_req,
      S_AXI_UFC_TX_TDATA  => aurora_ufc_tx_tdata,
      UFC_TX_MS           => aurora_ufc_tx_ms,
      S_AXI_UFC_TX_TVALID => aurora_ufc_tx_tvalid,
      S_AXI_UFC_TX_TREADY => aurora_ufc_tx_tready,
      -- UFC RX
      M_AXI_UFC_RX_TDATA  => aurora_ufc_rx_tdata,
      M_AXI_UFC_RX_TKEEP  => aurora_ufc_rx_tkeep,
      M_AXI_UFC_RX_TLAST  => aurora_ufc_rx_tlast,
      M_AXI_UFC_RX_TVALID => aurora_ufc_rx_tvalid,
      UFC_IN_PROGRESSn    => aurora_ufc_in_progress_n,
      -- GTX pins
      RXP                 => SMA_MGT_RX_P,
      RXN                 => SMA_MGT_RX_N,
      TXP                 => SMA_MGT_TX_P,
      TXN                 => SMA_MGT_TX_N,
      -- Status
      STATUS              => aurora_status
    );
  aurora_reset <= reset OR pulse_reg(15);
  fifo_over_ufc_inst : fifo_over_ufc
    PORT MAP (
      RESET            => aurora_reset,
      AURORA_USER_CLK  => aurora_user_clk,
      AURORA_TX_REQ    => aurora_ufc_tx_req,
      AURORA_TX_MS     => aurora_ufc_tx_ms,
      AURORA_TX_TREADY => aurora_ufc_tx_tready,
      AURORA_TX_TDATA  => aurora_ufc_tx_tdata,
      AURORA_TX_TVALID => aurora_ufc_tx_tvalid,
      AURORA_RX_TDATA  => aurora_ufc_rx_tdata,
      AURORA_RX_TVALID => aurora_ufc_rx_tvalid,
      FIFO_CLK         => control_fifo_rdclk,
      TX_FIFO_Q        => aurora_ufc_tx_fifo_q,
      TX_FIFO_WREN     => aurora_ufc_tx_fifo_wren,
      TX_FIFO_FULL     => aurora_ufc_tx_fifo_full,
      RX_FIFO_Q        => control_fifo_q(31 DOWNTO 0),
      RX_FIFO_RDEN     => control_fifo_rdreq,
      RX_FIFO_EMPTY    => control_fifo_empty,
      ERR              => OPEN -- LED8Bit(1)
    );
  fifo_over_ufc_tx_fifo : fifo36x512
    PORT MAP (
      rst    => aurora_reset,
      wr_clk => control_fifo_rdclk,
      rd_clk => control_clk,
      din    => x"0" & aurora_ufc_tx_fifo_q,
      wr_en  => aurora_ufc_tx_fifo_wren,
      rd_en  => cmd_fifo_rdreq,
      dout   => cmd_fifo_q,
      full   => aurora_ufc_tx_fifo_full,
      empty  => cmd_fifo_empty
    );

  -- -- debug
  -- aurora_ufc_tx_req <= pulse_reg(8);
  -- ufc_tx_tvalid_edge_sync_inst : edge_sync
  --   GENERIC MAP (
  --     EDGE => '0'
  --   )
  --   PORT MAP (
  --     RESET => reset,
  --     CLK   => aurora_user_clk,
  --     EI    => aurora_ufc_tx_req,
  --     SO    => aurora_ufc_tx_tvalid
  --   );
  -- aurora_ufc_tx_tdata <= x"0000_0000_0000" & config_reg(30*16+15 DOWNTO 30*16);
  -- aurora_ufc_tx_ms    <= config_reg(29*16+7 DOWNTO 29*16);  -- don't reverse bit-order here
  --
  dbg_ila1_inst : dbg_ila1
    PORT MAP (
      CLK    => clk_200MHz, -- aurora_user_clk,
      PROBE0 => dbg_ila1_probe0,
      PROBE1 => dbg_ila1_probe1
    );
  -- dbg_ila1_probe0 <=
  --   "00000" & aurora_status(2) & aurora_status(1) & aurora_status(0)
  --   & aurora_reset & aurora_ufc_in_progress_n & aurora_ufc_rx_tlast & aurora_ufc_rx_tvalid
  --   & aurora_ufc_tx_req & aurora_ufc_tx_tready & aurora_ufc_tx_tvalid & aurora_tx_tready;
  -- dbg_ila1_probe1 <= aurora_ufc_rx_tdata(7 DOWNTO 0) & aurora_ufc_tx_tdata(7 DOWNTO 0);
  ---------------------------------------------> gtx / aurora
  ---------------------------------------------< I2C
  i2c_sda_iobuf_inst : IOBUF
    GENERIC MAP(
      DRIVE      => 12,
      SLEW       => "SLOW"
    )
    PORT MAP(
      O  => i2c_sda_in,
      IO => I2C_SDA,
      I  => i2c_sda_out,
      T  => i2c_sda_t
    );
  i2c_scl_iobuf_inst : IOBUF
    GENERIC MAP(
      DRIVE      => 12,
      SLEW       => "SLOW"
    )
    PORT MAP(
      O  => OPEN,
      IO => I2C_SCL,
      I  => i2c_scl_out,
      T  => '0'
    );
  -- External clock IC
  si5338_clk_div_inst : clk_div
    GENERIC MAP (
      WIDTH => 32,
      PBITS => 8
    )
    PORT MAP (
      RESET   => reset,
      CLK     => clk156p25,
      DIV     => x"1b",
      CLK_DIV => LED8Bit(0)
    );
  -- Temperature and voltage sensors
  i2c1_sda_iobuf_inst : IOBUF
    GENERIC MAP(
      DRIVE      => 12,
      SLEW       => "SLOW"
    )
    PORT MAP(
      O  => i2c1_sda_in,
      IO => B14_L_P(19),
      I  => i2c1_sda_out,
      T  => i2c1_sda_t
    );
  i2c1_scl_iobuf_inst : IOBUF
    GENERIC MAP(
      DRIVE      => 12,
      SLEW       => "SLOW"
    )
    PORT MAP(
      O  => OPEN,
      IO => B14_L_P(14),
      I  => i2c1_scl_out,
      T  => '0'
    );
  i2c1_master_inst : i2c_master
    GENERIC MAP (
      INPUT_CLK_FREQENCY => 100_000_000,
      BUS_CLK_FREQUENCY  => 100_000
    )
    PORT MAP (
      CLK       => control_clk,
      RESET     => reset,
      START     => pulse_reg(2),
      MODE      => config_reg(16*2+1  DOWNTO 16*2),
      SL_RW     => config_reg(16*3+15),
      SL_ADDR   => config_reg(16*3+14 DOWNTO 16*3+8),
      REG_ADDR  => config_reg(16*3+7  DOWNTO 16*3),
      WR_DATA0  => config_reg(16*4+15 DOWNTO 16*4+8),
      WR_DATA1  => config_reg(16*4+7  DOWNTO 16*4),
      RD_DATA0  => status_reg(16*0+15 DOWNTO 16*0+8),
      RD_DATA1  => status_reg(16*0+7  DOWNTO 16*0),
      BUSY      => OPEN,
      ACK_ERROR => OPEN,
      SDA_in    => i2c1_sda_in,
      SDA_out   => i2c1_sda_out,
      SDA_t     => i2c1_sda_t,
      SCL       => i2c1_scl_out
    );
  ---------------------------------------------> I2C
  ---------------------------------------------< shiftreg driver for DAC8568
  B14_L_P(21) <= dac_din;
  B14_L_P(20) <= dac_sclk;
  B14_L_N(23) <= dac_sync_n;
  dac_din     <= spi_dout;
  dac_sclk    <= spi_sclk;
  dac_sync_n  <= spi_sync_n;
  dac8568_inst : fifo2shiftreg
    GENERIC MAP (
      DATA_WIDTH        => 32,          -- parallel data width
      CLK_DIV_WIDTH     => 16,
      DELAY_AFTER_SYNCn => 0,  -- number of SCLK cycles' wait after falling edge OF SYNCn
      SCLK_IDLE_LEVEL   => '0',  -- High or Low for SCLK when not switching
      DOUT_DRIVE_EDGE   => '1',  -- 1/0 rising/falling edge of SCLK drives new DOUT bit
      DIN_CAPTURE_EDGE  => '0'  -- 1/0 rising/falling edge of SCLK captures new DIN bit
    )
    PORT MAP (
      CLK      => control_clk,          -- clock
      RESET    => reset,                -- reset
      -- input data interface
      WR_CLK   => control_clk,          -- FIFO write clock
      DINFIFO  => config_reg(16*1+15 DOWNTO 16*1),
      WR_EN    => '0',
      WR_PULSE => pulse_reg(1),  -- one pulse writes one word, regardless of pulse duration
      FULL     => OPEN,
      -- captured data
      BUSY     => OPEN,
      DATAOUT  => OPEN,
      -- serial interface
      CLK_DIV  => x"0006",
      SCLK     => spi_sclk,
      DOUT     => spi_dout,
      SYNCn    => spi_sync_n,
      DIN      => spi_din
    );
  ---------------------------------------------> shiftreg driver for DAC8568
  ---------------------------------------------< TMS serial io
  B14_L_N(4)  <= tms_pwr_on;
  B14_L_P(4)  <= tms_sio_a(2);
  B14_L_N(13) <= tms_sio_a(1);
  B14_L_P(13) <= tms_sio_a(0);
  B14_L_P(23) <= tms_sdi;
  tms_sdo     <= B14_L_N(19);
  B14_L_P(0)  <= tms_sck;
  tms_pwr_on  <= config_reg(16*0+0);
  tms_sio_a   <= config_reg(16*13+8+tms_sio_a'length-1 DOWNTO 16*13+8);
  tms_sio_drive_inst : shiftreg_drive
    GENERIC MAP (
      DATA_WIDTH        => 130,         -- parallel data width
      CLK_DIV_WIDTH     => 16,
      DELAY_AFTER_SYNCn => 0,  -- number of SCLK cycles' wait after falling edge OF SYNCn
      SCLK_IDLE_LEVEL   => '1',  -- High or Low for SCLK when not switching
      DOUT_DRIVE_EDGE   => '0',  -- 1/0 rising/falling edge of SCLK drives new DOUT bit
      DIN_CAPTURE_EDGE  => '1'  -- 1/0 rising/falling edge of SCLK captures new DIN bit
    )
    PORT MAP (
      CLK     => control_clk,           -- clock
      RESET   => reset,                 -- reset
      -- internal data interface
      CLK_DIV => x"00" & "00" & config_reg(16*13+7 DOWNTO 16*13+2),  -- SCLK freq is CLK / 2**(CLK_DIV)
      DATAIN  => config_reg(16*13+1 DOWNTO 16*5),
      START   => pulse_reg(3),
      BUSY    => status_reg(16*9+2),
      DATAOUT => status_reg(16*9+1 DOWNTO 16*1),
      -- external serial interface
      SCLK    => tms_sck,
      DOUT    => tms_sdi,
      SYNCn   => OPEN,
      DIN     => tms_sdo
    );
  ---------------------------------------------> TMS serial io
  ---------------------------------------------< TMS
  -- TMS reset, also function as serial io load
  tms_reset_obufds_inst : OBUFDS
    GENERIC MAP(
      IOSTANDARD => "DEFAULT",
      SLEW       => "SLOW"
    )
    PORT MAP (
      O  => B13_L_P(3),
      OB => B13_L_N(3),
      I  => tms_reset
    );
  tms_reset_width_pulse_sync_inst : width_pulse_sync
    GENERIC MAP (
      DATA_WIDTH => 8,
      MODE       => 0
    )
    PORT MAP (
      RESET => reset,
      CLK   => control_clk,
      PW    => x"ff",
      START => pulse_reg(0),
      BUSY  => OPEN,
      CLKO  => control_clk,
      RSTO  => OPEN,
      PO    => tms_reset
    );
  -- TMS SDM
  B12_L_P(0)          <= tms_sdm_clk_src_sel;
  tms_sdm_clk_src_sel <= config_reg(16*0+1);
  tms_sdm_clkff_div   <= config_reg(16*0+11 DOWNTO 16*0+8);
  tms_sdm_recv_inst : tms_sdm_recv
    GENERIC MAP (
      NCH => 19
    )
    PORT MAP (
      RESET         => reset,
      CLK           => control_clk,  -- DELAY_* must be synchronous to this clock
      REFCLK        => clk_200MHz,   -- REFCLK (200MHz) for IDELAYCTRL
      DELAY_CHANNEL => config_reg(16*14+15 DOWNTO 16*14+8), -- input iodelay channel selection
      DELAY_VALUE   => config_reg(16*14+4 DOWNTO 16*14),    -- input iodelay value
      DELAY_UPDATE  => pulse_reg(4),    -- a pulse to update the delay value
      CLKFF_DIV     => tms_sdm_clkff_div,
      CLKFF_P       => B12_L_P(16),
      CLKFF_N       => B12_L_N(16),
      CLK_LPBK_P    => B12_L_P(12),
      CLK_LPBK_N    => B12_L_N(12),
      CLK_LPBK      => tms_sdm_clk_lpbk,
      SDM_OUT1_P    => tms_sdm_out1_p,
      SDM_OUT1_N    => tms_sdm_out1_n,
      SDM_OUT2_P    => tms_sdm_out2_p,
      SDM_OUT2_N    => tms_sdm_out2_n,
      DOUT          => tms_sdm_out
    );
  tms_sdm_out1_p <= (
    0  => B12_L_P(18),
    1  => B12_L_P(9),
    2  => B12_L_P(20),
    3  => B13_L_P(23),
    4  => B13_L_P(21),
    5  => B13_L_P(12),
    6  => B12_L_P(5),
    7  => B12_L_P(7),
    8  => B12_L_P(21),
    9  => B12_L_P(24),
    10 => B13_L_P(6),
    11 => B13_L_P(9),
    12 => B13_L_P(16),
    13 => B13_L_P(22),
    14 => B13_L_P(10),
    15 => B13_L_P(8),
    16 => B13_L_P(4),
    17 => B12_L_P(11),
    18 => B12_L_P(13)
  );
  tms_sdm_out1_n <= (
    0  => B12_L_N(18),
    1  => B12_L_N(9),
    2  => B12_L_N(20),
    3  => B13_L_N(23),
    4  => B13_L_N(21),
    5  => B13_L_N(12),
    6  => B12_L_N(5),
    7  => B12_L_N(7),
    8  => B12_L_N(21),
    9  => B12_L_N(24),
    10 => B13_L_N(6),
    11 => B13_L_N(9),
    12 => B13_L_N(16),
    13 => B13_L_N(22),
    14 => B13_L_N(10),
    15 => B13_L_N(8),
    16 => B13_L_N(4),
    17 => B12_L_N(11),
    18 => B12_L_N(13)
  );
  tms_sdm_out2_p <= (
    0  => B12_L_P(17),
    1  => B12_L_P(8),
    2  => B12_L_P(22),
    3  => B13_L_P(13),
    4  => B13_L_P(11),
    5  => B13_L_P(15),
    6  => B12_L_P(3),
    7  => B12_L_P(10),
    8  => B12_L_P(23),
    9  => B12_L_P(19),
    10 => B13_L_P(17),
    11 => B13_L_P(18),
    12 => B13_L_P(14),
    13 => B13_L_P(24),
    14 => B13_L_P(7),
    15 => B13_L_P(20),
    16 => B13_L_P(2),
    17 => B12_L_P(2),
    18 => B12_L_P(14)
  );
  tms_sdm_out2_n <= (
    0  => B12_L_N(17),
    1  => B12_L_N(8),
    2  => B12_L_N(22),
    3  => B13_L_N(13),
    4  => B13_L_N(11),
    5  => B13_L_N(15),
    6  => B12_L_N(3),
    7  => B12_L_N(10),
    8  => B12_L_N(23),
    9  => B12_L_N(19),
    10 => B13_L_N(17),
    11 => B13_L_N(18),
    12 => B13_L_N(14),
    13 => B13_L_N(24),
    14 => B13_L_N(7),
    15 => B13_L_N(20),
    16 => B13_L_N(2),
    17 => B12_L_N(2),
    18 => B12_L_N(14)
  );
  -- ADC, external, LTC2325-16
  B16_L_N(6)    <= adc_clk_src_sel;
  B16_L_N(19)   <= adc_clk_src_sel;
  B12_L_P(25)   <= adc_sdrn_ddr;
  adc_clk_src_sel <= config_reg(16*0+2);
  adc_sdrn_ddr    <= config_reg(16*0+3);
  adc_clkff_div   <= config_reg(16*0+15 DOWNTO 16*0+12);
  adc_cnv_sipo_inst : adc_cnv_sipo
    GENERIC MAP (
      NCH => 20
    )
    PORT MAP (
      RESET         => reset,
      CLK           => control_clk,  -- DELAY_* must be synchronous to this clock
      REFCLK        => clk_200MHz,   -- REFCLK (200MHz) for IDELAYCTRL
      DELAY_CHANNEL => config_reg(16*14+15 DOWNTO 16*14+8), -- ADC data input iodelay channel selection
      DELAY_VALUE   => config_reg(16*14+4 DOWNTO 16*14),    -- ADC data input iodelay value
      DELAY_UPDATE  => pulse_reg(5),    -- a pulse to update the delay value
      CLKFF_DIV     => adc_clkff_div,
      CLKFF_P       => B16_L_P(13),
      CLKFF_N       => B16_L_N(13),
      CLK_LPBK_P    => B16_L_P(12),
      CLK_LPBK_N    => B16_L_N(12),
      CLK_LPBK      => adc_clk0_lpbk,
      CNV_N_P       => B16_L_P(17),
      CNV_N_N       => B16_L_N(17),
      CNV_N         => adc_cnv_n,
      INPUTS_P      => adc_sdo_p,
      INPUTS_N      => adc_sdo_n,
      INPUTS_OUT    => adc_sdo,
      DOUT          => adc_dout,
      DOUT_VALID    => adc_dout_valid
    );
  adc_sdo_p <= (
    0  => B12_L_P(4),
    1  => B12_L_P(1),
    2  => B12_L_P(6),
    3  => B15_L_P(23),
    4  => B12_L_P(15),
    5  => B15_L_P(21),
    6  => B15_L_P(14),
    7  => B15_L_P(12),
    8  => B15_L_P(13),
    9  => B15_L_P(11),
    10 => B15_L_P(5),
    11 => B15_L_P(20),
    12 => B16_L_P(18),
    13 => B15_L_P(7),
    14 => B16_L_P(14),
    15 => B16_L_P(23),
    16 => B16_L_P(11),
    17 => B16_L_P(21),
    18 => B13_L_P(5),
    19 => B13_L_P(1)
  );
  adc_sdo_n <= (
    0  => B12_L_N(4),
    1  => B12_L_N(1),
    2  => B12_L_N(6),
    3  => B15_L_N(23),
    4  => B12_L_N(15),
    5  => B15_L_N(21),
    6  => B15_L_N(14),
    7  => B15_L_N(12),
    8  => B15_L_N(13),
    9  => B15_L_N(11),
    10 => B15_L_N(5),
    11 => B15_L_N(20),
    12 => B16_L_N(18),
    13 => B15_L_N(7),
    14 => B16_L_N(14),
    15 => B16_L_N(23),
    16 => B16_L_N(11),
    17 => B16_L_N(21),
    18 => B13_L_N(5),
    19 => B13_L_N(1)
  );
  --
  dbg_ila1_probe0 <= adc_dout(16*19+15 DOWNTO 16*19);
  dbg_ila1_probe1 <= tms_sdm_out(5 DOWNTO 0) & tms_sdm_clk_lpbk & tms_sck
                     & i2c1_sda_in & i2c1_sda_out & i2c1_scl_out & adc_dout_valid
                     & adc_cnv_n & adc_clk0_lpbk & adc_sdo(19) & adc_sdo(0);
  ---------------------------------------------> TMS

  -- clock output
  refout_clk_div_inst : clk_div
    PORT MAP (
      RESET   => reset,
      CLK     => idata_adc_data_clk,
      DIV     => config_reg(16*15+3 DOWNTO 16*15),
      CLK_DIV => idata_adc_refout_clkdiv
    );
  clk_fwd_inst : clk_fwd                -- idata_adc_refout_clkdiv
    PORT MAP (R => reset, I => clk156p25, O => OPEN);
  clk_fwd_inst1 : clk_fwd GENERIC MAP (INV => true)
    PORT MAP (R => reset, I => clk156p25, O => OPEN);
  clk_fwd_inst2 : clk_fwd GENERIC MAP (INV => true)
    PORT MAP (R => reset, I => idata_adc_data_clk, O => OPEN);

  -- capture the rising edge of trigger
  trig_edge_sync_inst : edge_sync
    PORT MAP (
      RESET => reset,
      CLK   => control_clk,
      EI    => idata_trig_in,
      SO    => idata_trig_synced
    );
  idata_trig_allow    <= config_reg(32*6+30);
  idata_data_wr_start <= pulse_reg(3) OR (idata_trig_synced AND idata_trig_allow
                                          AND (NOT idata_data_wr_busy)
                                          AND (NOT idata_data_wr_wrapped));

  --led_obufs : FOR i IN 0 TO 7 GENERATE
  --  led_obuf : OBUF
  --    PORT MAP (
  --      I => usr_data_output(i),
  --      O => LED8Bit(i)
  --    );
  --END GENERATE led_obufs;
  --LED8Bit(5 DOWNTO 1) <= (OTHERS => '0');

END Behavioral;
